// qsys_top.v

// Generated using ACDS version 23.4 79

`timescale 1 ps / 1 ps
module qsys_top (
		output wire        wd_reset_reset_n,         //             wd_reset.reset_n
		output wire        hps_io_EMAC0_TX_CLK,      //               hps_io.EMAC0_TX_CLK
		output wire        hps_io_EMAC0_TXD0,        //                     .EMAC0_TXD0
		output wire        hps_io_EMAC0_TXD1,        //                     .EMAC0_TXD1
		output wire        hps_io_EMAC0_TXD2,        //                     .EMAC0_TXD2
		output wire        hps_io_EMAC0_TXD3,        //                     .EMAC0_TXD3
		input  wire        hps_io_EMAC0_RX_CTL,      //                     .EMAC0_RX_CTL
		output wire        hps_io_EMAC0_TX_CTL,      //                     .EMAC0_TX_CTL
		input  wire        hps_io_EMAC0_RX_CLK,      //                     .EMAC0_RX_CLK
		input  wire        hps_io_EMAC0_RXD0,        //                     .EMAC0_RXD0
		input  wire        hps_io_EMAC0_RXD1,        //                     .EMAC0_RXD1
		input  wire        hps_io_EMAC0_RXD2,        //                     .EMAC0_RXD2
		input  wire        hps_io_EMAC0_RXD3,        //                     .EMAC0_RXD3
		inout  wire        hps_io_EMAC0_MDIO,        //                     .EMAC0_MDIO
		output wire        hps_io_EMAC0_MDC,         //                     .EMAC0_MDC
		inout  wire        hps_io_SDMMC_CMD,         //                     .SDMMC_CMD
		inout  wire        hps_io_SDMMC_D0,          //                     .SDMMC_D0
		inout  wire        hps_io_SDMMC_D1,          //                     .SDMMC_D1
		inout  wire        hps_io_SDMMC_D2,          //                     .SDMMC_D2
		inout  wire        hps_io_SDMMC_D3,          //                     .SDMMC_D3
		output wire        hps_io_SDMMC_CCLK,        //                     .SDMMC_CCLK
		inout  wire        hps_io_USB0_DATA0,        //                     .USB0_DATA0
		inout  wire        hps_io_USB0_DATA1,        //                     .USB0_DATA1
		inout  wire        hps_io_USB0_DATA2,        //                     .USB0_DATA2
		inout  wire        hps_io_USB0_DATA3,        //                     .USB0_DATA3
		inout  wire        hps_io_USB0_DATA4,        //                     .USB0_DATA4
		inout  wire        hps_io_USB0_DATA5,        //                     .USB0_DATA5
		inout  wire        hps_io_USB0_DATA6,        //                     .USB0_DATA6
		inout  wire        hps_io_USB0_DATA7,        //                     .USB0_DATA7
		input  wire        hps_io_USB0_CLK,          //                     .USB0_CLK
		output wire        hps_io_USB0_STP,          //                     .USB0_STP
		input  wire        hps_io_USB0_DIR,          //                     .USB0_DIR
		input  wire        hps_io_USB0_NXT,          //                     .USB0_NXT
		input  wire        hps_io_UART0_RX,          //                     .UART0_RX
		output wire        hps_io_UART0_TX,          //                     .UART0_TX
		inout  wire        hps_io_I2C1_SDA,          //                     .I2C1_SDA
		inout  wire        hps_io_I2C1_SCL,          //                     .I2C1_SCL
		inout  wire        hps_io_gpio1_io0,         //                     .gpio1_io0
		inout  wire        hps_io_gpio1_io1,         //                     .gpio1_io1
		inout  wire        hps_io_gpio1_io4,         //                     .gpio1_io4
		inout  wire        hps_io_gpio1_io5,         //                     .gpio1_io5
		input  wire        hps_io_jtag_tck,          //                     .jtag_tck
		input  wire        hps_io_jtag_tms,          //                     .jtag_tms
		output wire        hps_io_jtag_tdo,          //                     .jtag_tdo
		input  wire        hps_io_jtag_tdi,          //                     .jtag_tdi
		input  wire        hps_io_hps_osc_clk,       //                     .hps_osc_clk
		inout  wire        hps_io_gpio1_io19,        //                     .gpio1_io19
		inout  wire        hps_io_gpio1_io20,        //                     .gpio1_io20
		inout  wire        hps_io_gpio1_io21,        //                     .gpio1_io21
		output wire        h2f_reset_reset,          //            h2f_reset.reset
		input  wire        clk_100_clk,              //              clk_100.clk
		input  wire        emif_hps_pll_ref_clk_clk, // emif_hps_pll_ref_clk.clk
		input  wire        emif_hps_oct_oct_rzqin,   //         emif_hps_oct.oct_rzqin
		output wire [0:0]  emif_hps_mem_mem_ck,      //         emif_hps_mem.mem_ck
		output wire [0:0]  emif_hps_mem_mem_ck_n,    //                     .mem_ck_n
		output wire [16:0] emif_hps_mem_mem_a,       //                     .mem_a
		output wire [0:0]  emif_hps_mem_mem_act_n,   //                     .mem_act_n
		output wire [1:0]  emif_hps_mem_mem_ba,      //                     .mem_ba
		output wire [0:0]  emif_hps_mem_mem_bg,      //                     .mem_bg
		output wire [0:0]  emif_hps_mem_mem_cke,     //                     .mem_cke
		output wire [0:0]  emif_hps_mem_mem_cs_n,    //                     .mem_cs_n
		output wire [0:0]  emif_hps_mem_mem_odt,     //                     .mem_odt
		output wire [0:0]  emif_hps_mem_mem_reset_n, //                     .mem_reset_n
		output wire [0:0]  emif_hps_mem_mem_par,     //                     .mem_par
		input  wire [0:0]  emif_hps_mem_mem_alert_n, //                     .mem_alert_n
		inout  wire [8:0]  emif_hps_mem_mem_dqs,     //                     .mem_dqs
		inout  wire [8:0]  emif_hps_mem_mem_dqs_n,   //                     .mem_dqs_n
		inout  wire [71:0] emif_hps_mem_mem_dq,      //                     .mem_dq
		inout  wire [8:0]  emif_hps_mem_mem_dbi_n,   //                     .mem_dbi_n
		output wire [3:0]  fpga_led_pio_export,      //         fpga_led_pio.export
		input  wire        reset_reset_n,            //                reset.reset_n
		output wire        ninit_done_ninit_done     //           ninit_done.ninit_done
	);

	wire           emif_calbus_0_emif_calbus_clk_clk;                // emif_calbus_0:calbus_clk -> emif_hps:calbus_clk
	wire           clk_100_out_clk_clk;                              // clk_100:out_clk -> [agilex_hps:f2h_axi_clk, agilex_hps:h2f_axi_clk, agilex_hps:h2f_lw_axi_clk, mm_interconnect_0:clk_100_out_clk_clk, mm_interconnect_1:clk_100_out_clk_clk, onchip_memory2_0:clk, pio_1:clk, rst_controller:clk, rst_in:clk]
	wire    [31:0] emif_calbus_0_emif_calbus_0_calbus_wdata;         // emif_calbus_0:calbus_wdata_0 -> emif_hps:calbus_wdata
	wire    [19:0] emif_calbus_0_emif_calbus_0_calbus_address;       // emif_calbus_0:calbus_address_0 -> emif_hps:calbus_address
	wire  [4095:0] emif_hps_emif_calbus_calbus_seq_param_tbl;        // emif_hps:calbus_seq_param_tbl -> emif_calbus_0:calbus_seq_param_tbl_0
	wire           emif_calbus_0_emif_calbus_0_calbus_read;          // emif_calbus_0:calbus_read_0 -> emif_hps:calbus_read
	wire           emif_calbus_0_emif_calbus_0_calbus_write;         // emif_calbus_0:calbus_write_0 -> emif_hps:calbus_write
	wire    [31:0] emif_hps_emif_calbus_calbus_rdata;                // emif_hps:calbus_rdata -> emif_calbus_0:calbus_rdata_0
	wire     [1:0] agilex_hps_hps_emif_gp_to_emif;                   // agilex_hps:hps_emif_gp_to_emif -> emif_hps:hps_to_emif_gp
	wire  [4095:0] emif_hps_hps_emif_emif_to_hps;                    // emif_hps:emif_to_hps -> agilex_hps:hps_emif_emif_to_hps
	wire     [0:0] emif_hps_hps_emif_emif_to_gp;                     // emif_hps:emif_to_hps_gp -> agilex_hps:hps_emif_emif_to_gp
	wire  [4095:0] agilex_hps_hps_emif_hps_to_emif;                  // agilex_hps:hps_emif_hps_to_emif -> emif_hps:hps_to_emif
	wire     [1:0] agilex_hps_h2f_axi_master_awburst;                // agilex_hps:h2f_AWBURST -> mm_interconnect_0:agilex_hps_h2f_axi_master_awburst
	wire     [7:0] agilex_hps_h2f_axi_master_arlen;                  // agilex_hps:h2f_ARLEN -> mm_interconnect_0:agilex_hps_h2f_axi_master_arlen
	wire     [3:0] agilex_hps_h2f_axi_master_wstrb;                  // agilex_hps:h2f_WSTRB -> mm_interconnect_0:agilex_hps_h2f_axi_master_wstrb
	wire           agilex_hps_h2f_axi_master_wready;                 // mm_interconnect_0:agilex_hps_h2f_axi_master_wready -> agilex_hps:h2f_WREADY
	wire     [3:0] agilex_hps_h2f_axi_master_rid;                    // mm_interconnect_0:agilex_hps_h2f_axi_master_rid -> agilex_hps:h2f_RID
	wire           agilex_hps_h2f_axi_master_rready;                 // agilex_hps:h2f_RREADY -> mm_interconnect_0:agilex_hps_h2f_axi_master_rready
	wire     [7:0] agilex_hps_h2f_axi_master_awlen;                  // agilex_hps:h2f_AWLEN -> mm_interconnect_0:agilex_hps_h2f_axi_master_awlen
	wire     [3:0] agilex_hps_h2f_axi_master_arcache;                // agilex_hps:h2f_ARCACHE -> mm_interconnect_0:agilex_hps_h2f_axi_master_arcache
	wire           agilex_hps_h2f_axi_master_wvalid;                 // agilex_hps:h2f_WVALID -> mm_interconnect_0:agilex_hps_h2f_axi_master_wvalid
	wire    [31:0] agilex_hps_h2f_axi_master_araddr;                 // agilex_hps:h2f_ARADDR -> mm_interconnect_0:agilex_hps_h2f_axi_master_araddr
	wire     [2:0] agilex_hps_h2f_axi_master_arprot;                 // agilex_hps:h2f_ARPROT -> mm_interconnect_0:agilex_hps_h2f_axi_master_arprot
	wire     [2:0] agilex_hps_h2f_axi_master_awprot;                 // agilex_hps:h2f_AWPROT -> mm_interconnect_0:agilex_hps_h2f_axi_master_awprot
	wire    [31:0] agilex_hps_h2f_axi_master_wdata;                  // agilex_hps:h2f_WDATA -> mm_interconnect_0:agilex_hps_h2f_axi_master_wdata
	wire           agilex_hps_h2f_axi_master_arvalid;                // agilex_hps:h2f_ARVALID -> mm_interconnect_0:agilex_hps_h2f_axi_master_arvalid
	wire     [3:0] agilex_hps_h2f_axi_master_awcache;                // agilex_hps:h2f_AWCACHE -> mm_interconnect_0:agilex_hps_h2f_axi_master_awcache
	wire     [3:0] agilex_hps_h2f_axi_master_arid;                   // agilex_hps:h2f_ARID -> mm_interconnect_0:agilex_hps_h2f_axi_master_arid
	wire           agilex_hps_h2f_axi_master_arlock;                 // agilex_hps:h2f_ARLOCK -> mm_interconnect_0:agilex_hps_h2f_axi_master_arlock
	wire           agilex_hps_h2f_axi_master_awlock;                 // agilex_hps:h2f_AWLOCK -> mm_interconnect_0:agilex_hps_h2f_axi_master_awlock
	wire    [31:0] agilex_hps_h2f_axi_master_awaddr;                 // agilex_hps:h2f_AWADDR -> mm_interconnect_0:agilex_hps_h2f_axi_master_awaddr
	wire     [1:0] agilex_hps_h2f_axi_master_bresp;                  // mm_interconnect_0:agilex_hps_h2f_axi_master_bresp -> agilex_hps:h2f_BRESP
	wire           agilex_hps_h2f_axi_master_arready;                // mm_interconnect_0:agilex_hps_h2f_axi_master_arready -> agilex_hps:h2f_ARREADY
	wire    [31:0] agilex_hps_h2f_axi_master_rdata;                  // mm_interconnect_0:agilex_hps_h2f_axi_master_rdata -> agilex_hps:h2f_RDATA
	wire           agilex_hps_h2f_axi_master_awready;                // mm_interconnect_0:agilex_hps_h2f_axi_master_awready -> agilex_hps:h2f_AWREADY
	wire     [1:0] agilex_hps_h2f_axi_master_arburst;                // agilex_hps:h2f_ARBURST -> mm_interconnect_0:agilex_hps_h2f_axi_master_arburst
	wire     [2:0] agilex_hps_h2f_axi_master_arsize;                 // agilex_hps:h2f_ARSIZE -> mm_interconnect_0:agilex_hps_h2f_axi_master_arsize
	wire           agilex_hps_h2f_axi_master_bready;                 // agilex_hps:h2f_BREADY -> mm_interconnect_0:agilex_hps_h2f_axi_master_bready
	wire           agilex_hps_h2f_axi_master_rlast;                  // mm_interconnect_0:agilex_hps_h2f_axi_master_rlast -> agilex_hps:h2f_RLAST
	wire           agilex_hps_h2f_axi_master_wlast;                  // agilex_hps:h2f_WLAST -> mm_interconnect_0:agilex_hps_h2f_axi_master_wlast
	wire     [1:0] agilex_hps_h2f_axi_master_rresp;                  // mm_interconnect_0:agilex_hps_h2f_axi_master_rresp -> agilex_hps:h2f_RRESP
	wire     [3:0] agilex_hps_h2f_axi_master_awid;                   // agilex_hps:h2f_AWID -> mm_interconnect_0:agilex_hps_h2f_axi_master_awid
	wire     [3:0] agilex_hps_h2f_axi_master_bid;                    // mm_interconnect_0:agilex_hps_h2f_axi_master_bid -> agilex_hps:h2f_BID
	wire           agilex_hps_h2f_axi_master_bvalid;                 // mm_interconnect_0:agilex_hps_h2f_axi_master_bvalid -> agilex_hps:h2f_BVALID
	wire     [2:0] agilex_hps_h2f_axi_master_awsize;                 // agilex_hps:h2f_AWSIZE -> mm_interconnect_0:agilex_hps_h2f_axi_master_awsize
	wire           agilex_hps_h2f_axi_master_awvalid;                // agilex_hps:h2f_AWVALID -> mm_interconnect_0:agilex_hps_h2f_axi_master_awvalid
	wire           agilex_hps_h2f_axi_master_rvalid;                 // mm_interconnect_0:agilex_hps_h2f_axi_master_rvalid -> agilex_hps:h2f_RVALID
	wire           mm_interconnect_0_onchip_memory2_0_s1_chipselect; // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire    [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;   // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire     [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;    // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire     [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable; // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire           mm_interconnect_0_onchip_memory2_0_s1_write;      // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire    [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;  // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire           mm_interconnect_0_onchip_memory2_0_s1_clken;      // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire           rst_in_out_reset_reset;                           // rst_in:out_reset_n -> [mm_interconnect_0:agilex_hps_h2f_axi_master_translator_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:agilex_hps_h2f_axi_reset_reset_bridge_in_reset_reset, mm_interconnect_1:agilex_hps_h2f_lw_axi_master_translator_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:agilex_hps_h2f_lw_axi_reset_reset_bridge_in_reset_reset, rst_controller:reset_in0]
	wire     [1:0] agilex_hps_h2f_lw_axi_master_awburst;             // agilex_hps:h2f_lw_AWBURST -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_awburst
	wire     [7:0] agilex_hps_h2f_lw_axi_master_arlen;               // agilex_hps:h2f_lw_ARLEN -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_arlen
	wire     [3:0] agilex_hps_h2f_lw_axi_master_wstrb;               // agilex_hps:h2f_lw_WSTRB -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_wstrb
	wire           agilex_hps_h2f_lw_axi_master_wready;              // mm_interconnect_1:agilex_hps_h2f_lw_axi_master_wready -> agilex_hps:h2f_lw_WREADY
	wire     [3:0] agilex_hps_h2f_lw_axi_master_rid;                 // mm_interconnect_1:agilex_hps_h2f_lw_axi_master_rid -> agilex_hps:h2f_lw_RID
	wire           agilex_hps_h2f_lw_axi_master_rready;              // agilex_hps:h2f_lw_RREADY -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_rready
	wire     [7:0] agilex_hps_h2f_lw_axi_master_awlen;               // agilex_hps:h2f_lw_AWLEN -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_awlen
	wire     [3:0] agilex_hps_h2f_lw_axi_master_arcache;             // agilex_hps:h2f_lw_ARCACHE -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_arcache
	wire           agilex_hps_h2f_lw_axi_master_wvalid;              // agilex_hps:h2f_lw_WVALID -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_wvalid
	wire    [20:0] agilex_hps_h2f_lw_axi_master_araddr;              // agilex_hps:h2f_lw_ARADDR -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_araddr
	wire     [2:0] agilex_hps_h2f_lw_axi_master_arprot;              // agilex_hps:h2f_lw_ARPROT -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_arprot
	wire     [2:0] agilex_hps_h2f_lw_axi_master_awprot;              // agilex_hps:h2f_lw_AWPROT -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_awprot
	wire    [31:0] agilex_hps_h2f_lw_axi_master_wdata;               // agilex_hps:h2f_lw_WDATA -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_wdata
	wire           agilex_hps_h2f_lw_axi_master_arvalid;             // agilex_hps:h2f_lw_ARVALID -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_arvalid
	wire     [3:0] agilex_hps_h2f_lw_axi_master_awcache;             // agilex_hps:h2f_lw_AWCACHE -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_awcache
	wire     [3:0] agilex_hps_h2f_lw_axi_master_arid;                // agilex_hps:h2f_lw_ARID -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_arid
	wire           agilex_hps_h2f_lw_axi_master_arlock;              // agilex_hps:h2f_lw_ARLOCK -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_arlock
	wire           agilex_hps_h2f_lw_axi_master_awlock;              // agilex_hps:h2f_lw_AWLOCK -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_awlock
	wire    [20:0] agilex_hps_h2f_lw_axi_master_awaddr;              // agilex_hps:h2f_lw_AWADDR -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_awaddr
	wire     [1:0] agilex_hps_h2f_lw_axi_master_bresp;               // mm_interconnect_1:agilex_hps_h2f_lw_axi_master_bresp -> agilex_hps:h2f_lw_BRESP
	wire           agilex_hps_h2f_lw_axi_master_arready;             // mm_interconnect_1:agilex_hps_h2f_lw_axi_master_arready -> agilex_hps:h2f_lw_ARREADY
	wire    [31:0] agilex_hps_h2f_lw_axi_master_rdata;               // mm_interconnect_1:agilex_hps_h2f_lw_axi_master_rdata -> agilex_hps:h2f_lw_RDATA
	wire           agilex_hps_h2f_lw_axi_master_awready;             // mm_interconnect_1:agilex_hps_h2f_lw_axi_master_awready -> agilex_hps:h2f_lw_AWREADY
	wire     [1:0] agilex_hps_h2f_lw_axi_master_arburst;             // agilex_hps:h2f_lw_ARBURST -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_arburst
	wire     [2:0] agilex_hps_h2f_lw_axi_master_arsize;              // agilex_hps:h2f_lw_ARSIZE -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_arsize
	wire           agilex_hps_h2f_lw_axi_master_bready;              // agilex_hps:h2f_lw_BREADY -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_bready
	wire           agilex_hps_h2f_lw_axi_master_rlast;               // mm_interconnect_1:agilex_hps_h2f_lw_axi_master_rlast -> agilex_hps:h2f_lw_RLAST
	wire           agilex_hps_h2f_lw_axi_master_wlast;               // agilex_hps:h2f_lw_WLAST -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_wlast
	wire     [1:0] agilex_hps_h2f_lw_axi_master_rresp;               // mm_interconnect_1:agilex_hps_h2f_lw_axi_master_rresp -> agilex_hps:h2f_lw_RRESP
	wire     [3:0] agilex_hps_h2f_lw_axi_master_awid;                // agilex_hps:h2f_lw_AWID -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_awid
	wire     [3:0] agilex_hps_h2f_lw_axi_master_bid;                 // mm_interconnect_1:agilex_hps_h2f_lw_axi_master_bid -> agilex_hps:h2f_lw_BID
	wire           agilex_hps_h2f_lw_axi_master_bvalid;              // mm_interconnect_1:agilex_hps_h2f_lw_axi_master_bvalid -> agilex_hps:h2f_lw_BVALID
	wire     [2:0] agilex_hps_h2f_lw_axi_master_awsize;              // agilex_hps:h2f_lw_AWSIZE -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_awsize
	wire           agilex_hps_h2f_lw_axi_master_awvalid;             // agilex_hps:h2f_lw_AWVALID -> mm_interconnect_1:agilex_hps_h2f_lw_axi_master_awvalid
	wire           agilex_hps_h2f_lw_axi_master_rvalid;              // mm_interconnect_1:agilex_hps_h2f_lw_axi_master_rvalid -> agilex_hps:h2f_lw_RVALID
	wire           mm_interconnect_1_pio_1_s1_chipselect;            // mm_interconnect_1:pio_1_s1_chipselect -> pio_1:chipselect
	wire    [31:0] mm_interconnect_1_pio_1_s1_readdata;              // pio_1:readdata -> mm_interconnect_1:pio_1_s1_readdata
	wire     [1:0] mm_interconnect_1_pio_1_s1_address;               // mm_interconnect_1:pio_1_s1_address -> pio_1:address
	wire           mm_interconnect_1_pio_1_s1_write;                 // mm_interconnect_1:pio_1_s1_write -> pio_1:write_n
	wire    [31:0] mm_interconnect_1_pio_1_s1_writedata;             // mm_interconnect_1:pio_1_s1_writedata -> pio_1:writedata
	wire           rst_controller_reset_out_reset;                   // rst_controller:reset_out -> [agilex_hps:f2h_axi_rst_n, agilex_hps:h2f_axi_rst_n, agilex_hps:h2f_lw_axi_rst_n, onchip_memory2_0:reset, pio_1:reset_n, rst_translator:in_reset]
	wire           rst_controller_reset_out_reset_req;               // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	agilex_hps agilex_hps (
		.h2f_watchdog_rst     (wd_reset_reset_n),                     //  output,     width = 1,  h2f_watchdog_rst.reset_n
		.hps_emif_emif_to_hps (emif_hps_hps_emif_emif_to_hps),        //   input,  width = 4096,          hps_emif.emif_to_hps
		.hps_emif_hps_to_emif (agilex_hps_hps_emif_hps_to_emif),      //  output,  width = 4096,                  .hps_to_emif
		.hps_emif_emif_to_gp  (emif_hps_hps_emif_emif_to_gp),         //   input,     width = 1,                  .emif_to_gp
		.hps_emif_gp_to_emif  (agilex_hps_hps_emif_gp_to_emif),       //  output,     width = 2,                  .gp_to_emif
		.EMAC0_TX_CLK         (hps_io_EMAC0_TX_CLK),                  //  output,     width = 1,            hps_io.EMAC0_TX_CLK
		.EMAC0_TXD0           (hps_io_EMAC0_TXD0),                    //  output,     width = 1,                  .EMAC0_TXD0
		.EMAC0_TXD1           (hps_io_EMAC0_TXD1),                    //  output,     width = 1,                  .EMAC0_TXD1
		.EMAC0_TXD2           (hps_io_EMAC0_TXD2),                    //  output,     width = 1,                  .EMAC0_TXD2
		.EMAC0_TXD3           (hps_io_EMAC0_TXD3),                    //  output,     width = 1,                  .EMAC0_TXD3
		.EMAC0_RX_CTL         (hps_io_EMAC0_RX_CTL),                  //   input,     width = 1,                  .EMAC0_RX_CTL
		.EMAC0_TX_CTL         (hps_io_EMAC0_TX_CTL),                  //  output,     width = 1,                  .EMAC0_TX_CTL
		.EMAC0_RX_CLK         (hps_io_EMAC0_RX_CLK),                  //   input,     width = 1,                  .EMAC0_RX_CLK
		.EMAC0_RXD0           (hps_io_EMAC0_RXD0),                    //   input,     width = 1,                  .EMAC0_RXD0
		.EMAC0_RXD1           (hps_io_EMAC0_RXD1),                    //   input,     width = 1,                  .EMAC0_RXD1
		.EMAC0_RXD2           (hps_io_EMAC0_RXD2),                    //   input,     width = 1,                  .EMAC0_RXD2
		.EMAC0_RXD3           (hps_io_EMAC0_RXD3),                    //   input,     width = 1,                  .EMAC0_RXD3
		.EMAC0_MDIO           (hps_io_EMAC0_MDIO),                    //   inout,     width = 1,                  .EMAC0_MDIO
		.EMAC0_MDC            (hps_io_EMAC0_MDC),                     //  output,     width = 1,                  .EMAC0_MDC
		.SDMMC_CMD            (hps_io_SDMMC_CMD),                     //   inout,     width = 1,                  .SDMMC_CMD
		.SDMMC_D0             (hps_io_SDMMC_D0),                      //   inout,     width = 1,                  .SDMMC_D0
		.SDMMC_D1             (hps_io_SDMMC_D1),                      //   inout,     width = 1,                  .SDMMC_D1
		.SDMMC_D2             (hps_io_SDMMC_D2),                      //   inout,     width = 1,                  .SDMMC_D2
		.SDMMC_D3             (hps_io_SDMMC_D3),                      //   inout,     width = 1,                  .SDMMC_D3
		.SDMMC_CCLK           (hps_io_SDMMC_CCLK),                    //  output,     width = 1,                  .SDMMC_CCLK
		.USB0_DATA0           (hps_io_USB0_DATA0),                    //   inout,     width = 1,                  .USB0_DATA0
		.USB0_DATA1           (hps_io_USB0_DATA1),                    //   inout,     width = 1,                  .USB0_DATA1
		.USB0_DATA2           (hps_io_USB0_DATA2),                    //   inout,     width = 1,                  .USB0_DATA2
		.USB0_DATA3           (hps_io_USB0_DATA3),                    //   inout,     width = 1,                  .USB0_DATA3
		.USB0_DATA4           (hps_io_USB0_DATA4),                    //   inout,     width = 1,                  .USB0_DATA4
		.USB0_DATA5           (hps_io_USB0_DATA5),                    //   inout,     width = 1,                  .USB0_DATA5
		.USB0_DATA6           (hps_io_USB0_DATA6),                    //   inout,     width = 1,                  .USB0_DATA6
		.USB0_DATA7           (hps_io_USB0_DATA7),                    //   inout,     width = 1,                  .USB0_DATA7
		.USB0_CLK             (hps_io_USB0_CLK),                      //   input,     width = 1,                  .USB0_CLK
		.USB0_STP             (hps_io_USB0_STP),                      //  output,     width = 1,                  .USB0_STP
		.USB0_DIR             (hps_io_USB0_DIR),                      //   input,     width = 1,                  .USB0_DIR
		.USB0_NXT             (hps_io_USB0_NXT),                      //   input,     width = 1,                  .USB0_NXT
		.UART0_RX             (hps_io_UART0_RX),                      //   input,     width = 1,                  .UART0_RX
		.UART0_TX             (hps_io_UART0_TX),                      //  output,     width = 1,                  .UART0_TX
		.I2C1_SDA             (hps_io_I2C1_SDA),                      //   inout,     width = 1,                  .I2C1_SDA
		.I2C1_SCL             (hps_io_I2C1_SCL),                      //   inout,     width = 1,                  .I2C1_SCL
		.gpio1_io0            (hps_io_gpio1_io0),                     //   inout,     width = 1,                  .gpio1_io0
		.gpio1_io1            (hps_io_gpio1_io1),                     //   inout,     width = 1,                  .gpio1_io1
		.gpio1_io4            (hps_io_gpio1_io4),                     //   inout,     width = 1,                  .gpio1_io4
		.gpio1_io5            (hps_io_gpio1_io5),                     //   inout,     width = 1,                  .gpio1_io5
		.jtag_tck             (hps_io_jtag_tck),                      //   input,     width = 1,                  .jtag_tck
		.jtag_tms             (hps_io_jtag_tms),                      //   input,     width = 1,                  .jtag_tms
		.jtag_tdo             (hps_io_jtag_tdo),                      //  output,     width = 1,                  .jtag_tdo
		.jtag_tdi             (hps_io_jtag_tdi),                      //   input,     width = 1,                  .jtag_tdi
		.hps_osc_clk          (hps_io_hps_osc_clk),                   //   input,     width = 1,                  .hps_osc_clk
		.gpio1_io19           (hps_io_gpio1_io19),                    //   inout,     width = 1,                  .gpio1_io19
		.gpio1_io20           (hps_io_gpio1_io20),                    //   inout,     width = 1,                  .gpio1_io20
		.gpio1_io21           (hps_io_gpio1_io21),                    //   inout,     width = 1,                  .gpio1_io21
		.h2f_rst              (h2f_reset_reset),                      //  output,     width = 1,         h2f_reset.reset
		.h2f_axi_clk          (clk_100_out_clk_clk),                  //   input,     width = 1,     h2f_axi_clock.clk
		.h2f_axi_rst_n        (~rst_controller_reset_out_reset),      //   input,     width = 1,     h2f_axi_reset.reset_n
		.h2f_AWID             (agilex_hps_h2f_axi_master_awid),       //  output,     width = 4,    h2f_axi_master.awid
		.h2f_AWADDR           (agilex_hps_h2f_axi_master_awaddr),     //  output,    width = 32,                  .awaddr
		.h2f_AWLEN            (agilex_hps_h2f_axi_master_awlen),      //  output,     width = 8,                  .awlen
		.h2f_AWSIZE           (agilex_hps_h2f_axi_master_awsize),     //  output,     width = 3,                  .awsize
		.h2f_AWBURST          (agilex_hps_h2f_axi_master_awburst),    //  output,     width = 2,                  .awburst
		.h2f_AWLOCK           (agilex_hps_h2f_axi_master_awlock),     //  output,     width = 1,                  .awlock
		.h2f_AWCACHE          (agilex_hps_h2f_axi_master_awcache),    //  output,     width = 4,                  .awcache
		.h2f_AWPROT           (agilex_hps_h2f_axi_master_awprot),     //  output,     width = 3,                  .awprot
		.h2f_AWVALID          (agilex_hps_h2f_axi_master_awvalid),    //  output,     width = 1,                  .awvalid
		.h2f_AWREADY          (agilex_hps_h2f_axi_master_awready),    //   input,     width = 1,                  .awready
		.h2f_WDATA            (agilex_hps_h2f_axi_master_wdata),      //  output,    width = 32,                  .wdata
		.h2f_WSTRB            (agilex_hps_h2f_axi_master_wstrb),      //  output,     width = 4,                  .wstrb
		.h2f_WLAST            (agilex_hps_h2f_axi_master_wlast),      //  output,     width = 1,                  .wlast
		.h2f_WVALID           (agilex_hps_h2f_axi_master_wvalid),     //  output,     width = 1,                  .wvalid
		.h2f_WREADY           (agilex_hps_h2f_axi_master_wready),     //   input,     width = 1,                  .wready
		.h2f_BID              (agilex_hps_h2f_axi_master_bid),        //   input,     width = 4,                  .bid
		.h2f_BRESP            (agilex_hps_h2f_axi_master_bresp),      //   input,     width = 2,                  .bresp
		.h2f_BVALID           (agilex_hps_h2f_axi_master_bvalid),     //   input,     width = 1,                  .bvalid
		.h2f_BREADY           (agilex_hps_h2f_axi_master_bready),     //  output,     width = 1,                  .bready
		.h2f_ARID             (agilex_hps_h2f_axi_master_arid),       //  output,     width = 4,                  .arid
		.h2f_ARADDR           (agilex_hps_h2f_axi_master_araddr),     //  output,    width = 32,                  .araddr
		.h2f_ARLEN            (agilex_hps_h2f_axi_master_arlen),      //  output,     width = 8,                  .arlen
		.h2f_ARSIZE           (agilex_hps_h2f_axi_master_arsize),     //  output,     width = 3,                  .arsize
		.h2f_ARBURST          (agilex_hps_h2f_axi_master_arburst),    //  output,     width = 2,                  .arburst
		.h2f_ARLOCK           (agilex_hps_h2f_axi_master_arlock),     //  output,     width = 1,                  .arlock
		.h2f_ARCACHE          (agilex_hps_h2f_axi_master_arcache),    //  output,     width = 4,                  .arcache
		.h2f_ARPROT           (agilex_hps_h2f_axi_master_arprot),     //  output,     width = 3,                  .arprot
		.h2f_ARVALID          (agilex_hps_h2f_axi_master_arvalid),    //  output,     width = 1,                  .arvalid
		.h2f_ARREADY          (agilex_hps_h2f_axi_master_arready),    //   input,     width = 1,                  .arready
		.h2f_RID              (agilex_hps_h2f_axi_master_rid),        //   input,     width = 4,                  .rid
		.h2f_RDATA            (agilex_hps_h2f_axi_master_rdata),      //   input,    width = 32,                  .rdata
		.h2f_RRESP            (agilex_hps_h2f_axi_master_rresp),      //   input,     width = 2,                  .rresp
		.h2f_RLAST            (agilex_hps_h2f_axi_master_rlast),      //   input,     width = 1,                  .rlast
		.h2f_RVALID           (agilex_hps_h2f_axi_master_rvalid),     //   input,     width = 1,                  .rvalid
		.h2f_RREADY           (agilex_hps_h2f_axi_master_rready),     //  output,     width = 1,                  .rready
		.h2f_lw_axi_clk       (clk_100_out_clk_clk),                  //   input,     width = 1,  h2f_lw_axi_clock.clk
		.h2f_lw_axi_rst_n     (~rst_controller_reset_out_reset),      //   input,     width = 1,  h2f_lw_axi_reset.reset_n
		.h2f_lw_AWID          (agilex_hps_h2f_lw_axi_master_awid),    //  output,     width = 4, h2f_lw_axi_master.awid
		.h2f_lw_AWADDR        (agilex_hps_h2f_lw_axi_master_awaddr),  //  output,    width = 21,                  .awaddr
		.h2f_lw_AWLEN         (agilex_hps_h2f_lw_axi_master_awlen),   //  output,     width = 8,                  .awlen
		.h2f_lw_AWSIZE        (agilex_hps_h2f_lw_axi_master_awsize),  //  output,     width = 3,                  .awsize
		.h2f_lw_AWBURST       (agilex_hps_h2f_lw_axi_master_awburst), //  output,     width = 2,                  .awburst
		.h2f_lw_AWLOCK        (agilex_hps_h2f_lw_axi_master_awlock),  //  output,     width = 1,                  .awlock
		.h2f_lw_AWCACHE       (agilex_hps_h2f_lw_axi_master_awcache), //  output,     width = 4,                  .awcache
		.h2f_lw_AWPROT        (agilex_hps_h2f_lw_axi_master_awprot),  //  output,     width = 3,                  .awprot
		.h2f_lw_AWVALID       (agilex_hps_h2f_lw_axi_master_awvalid), //  output,     width = 1,                  .awvalid
		.h2f_lw_AWREADY       (agilex_hps_h2f_lw_axi_master_awready), //   input,     width = 1,                  .awready
		.h2f_lw_WDATA         (agilex_hps_h2f_lw_axi_master_wdata),   //  output,    width = 32,                  .wdata
		.h2f_lw_WSTRB         (agilex_hps_h2f_lw_axi_master_wstrb),   //  output,     width = 4,                  .wstrb
		.h2f_lw_WLAST         (agilex_hps_h2f_lw_axi_master_wlast),   //  output,     width = 1,                  .wlast
		.h2f_lw_WVALID        (agilex_hps_h2f_lw_axi_master_wvalid),  //  output,     width = 1,                  .wvalid
		.h2f_lw_WREADY        (agilex_hps_h2f_lw_axi_master_wready),  //   input,     width = 1,                  .wready
		.h2f_lw_BID           (agilex_hps_h2f_lw_axi_master_bid),     //   input,     width = 4,                  .bid
		.h2f_lw_BRESP         (agilex_hps_h2f_lw_axi_master_bresp),   //   input,     width = 2,                  .bresp
		.h2f_lw_BVALID        (agilex_hps_h2f_lw_axi_master_bvalid),  //   input,     width = 1,                  .bvalid
		.h2f_lw_BREADY        (agilex_hps_h2f_lw_axi_master_bready),  //  output,     width = 1,                  .bready
		.h2f_lw_ARID          (agilex_hps_h2f_lw_axi_master_arid),    //  output,     width = 4,                  .arid
		.h2f_lw_ARADDR        (agilex_hps_h2f_lw_axi_master_araddr),  //  output,    width = 21,                  .araddr
		.h2f_lw_ARLEN         (agilex_hps_h2f_lw_axi_master_arlen),   //  output,     width = 8,                  .arlen
		.h2f_lw_ARSIZE        (agilex_hps_h2f_lw_axi_master_arsize),  //  output,     width = 3,                  .arsize
		.h2f_lw_ARBURST       (agilex_hps_h2f_lw_axi_master_arburst), //  output,     width = 2,                  .arburst
		.h2f_lw_ARLOCK        (agilex_hps_h2f_lw_axi_master_arlock),  //  output,     width = 1,                  .arlock
		.h2f_lw_ARCACHE       (agilex_hps_h2f_lw_axi_master_arcache), //  output,     width = 4,                  .arcache
		.h2f_lw_ARPROT        (agilex_hps_h2f_lw_axi_master_arprot),  //  output,     width = 3,                  .arprot
		.h2f_lw_ARVALID       (agilex_hps_h2f_lw_axi_master_arvalid), //  output,     width = 1,                  .arvalid
		.h2f_lw_ARREADY       (agilex_hps_h2f_lw_axi_master_arready), //   input,     width = 1,                  .arready
		.h2f_lw_RID           (agilex_hps_h2f_lw_axi_master_rid),     //   input,     width = 4,                  .rid
		.h2f_lw_RDATA         (agilex_hps_h2f_lw_axi_master_rdata),   //   input,    width = 32,                  .rdata
		.h2f_lw_RRESP         (agilex_hps_h2f_lw_axi_master_rresp),   //   input,     width = 2,                  .rresp
		.h2f_lw_RLAST         (agilex_hps_h2f_lw_axi_master_rlast),   //   input,     width = 1,                  .rlast
		.h2f_lw_RVALID        (agilex_hps_h2f_lw_axi_master_rvalid),  //   input,     width = 1,                  .rvalid
		.h2f_lw_RREADY        (agilex_hps_h2f_lw_axi_master_rready),  //  output,     width = 1,                  .rready
		.f2h_axi_clk          (clk_100_out_clk_clk),                  //   input,     width = 1,     f2h_axi_clock.clk
		.f2h_axi_rst_n        (~rst_controller_reset_out_reset),      //   input,     width = 1,     f2h_axi_reset.reset_n
		.f2h_AWID             (),                                     //   input,     width = 5,     f2h_axi_slave.awid
		.f2h_AWADDR           (),                                     //   input,    width = 32,                  .awaddr
		.f2h_AWLEN            (),                                     //   input,     width = 8,                  .awlen
		.f2h_AWSIZE           (),                                     //   input,     width = 3,                  .awsize
		.f2h_AWBURST          (),                                     //   input,     width = 2,                  .awburst
		.f2h_AWLOCK           (),                                     //   input,     width = 1,                  .awlock
		.f2h_AWCACHE          (),                                     //   input,     width = 4,                  .awcache
		.f2h_AWPROT           (),                                     //   input,     width = 3,                  .awprot
		.f2h_AWVALID          (),                                     //   input,     width = 1,                  .awvalid
		.f2h_AWREADY          (),                                     //  output,     width = 1,                  .awready
		.f2h_AWQOS            (),                                     //   input,     width = 4,                  .awqos
		.f2h_WDATA            (),                                     //   input,   width = 128,                  .wdata
		.f2h_WSTRB            (),                                     //   input,    width = 16,                  .wstrb
		.f2h_WLAST            (),                                     //   input,     width = 1,                  .wlast
		.f2h_WVALID           (),                                     //   input,     width = 1,                  .wvalid
		.f2h_WREADY           (),                                     //  output,     width = 1,                  .wready
		.f2h_BID              (),                                     //  output,     width = 5,                  .bid
		.f2h_BRESP            (),                                     //  output,     width = 2,                  .bresp
		.f2h_BVALID           (),                                     //  output,     width = 1,                  .bvalid
		.f2h_BREADY           (),                                     //   input,     width = 1,                  .bready
		.f2h_ARID             (),                                     //   input,     width = 5,                  .arid
		.f2h_ARADDR           (),                                     //   input,    width = 32,                  .araddr
		.f2h_ARLEN            (),                                     //   input,     width = 8,                  .arlen
		.f2h_ARSIZE           (),                                     //   input,     width = 3,                  .arsize
		.f2h_ARBURST          (),                                     //   input,     width = 2,                  .arburst
		.f2h_ARLOCK           (),                                     //   input,     width = 1,                  .arlock
		.f2h_ARCACHE          (),                                     //   input,     width = 4,                  .arcache
		.f2h_ARPROT           (),                                     //   input,     width = 3,                  .arprot
		.f2h_ARVALID          (),                                     //   input,     width = 1,                  .arvalid
		.f2h_ARREADY          (),                                     //  output,     width = 1,                  .arready
		.f2h_ARQOS            (),                                     //   input,     width = 4,                  .arqos
		.f2h_RID              (),                                     //  output,     width = 5,                  .rid
		.f2h_RDATA            (),                                     //  output,   width = 128,                  .rdata
		.f2h_RRESP            (),                                     //  output,     width = 2,                  .rresp
		.f2h_RLAST            (),                                     //  output,     width = 1,                  .rlast
		.f2h_RVALID           (),                                     //  output,     width = 1,                  .rvalid
		.f2h_RREADY           (),                                     //   input,     width = 1,                  .rready
		.f2h_ARUSER           (),                                     //   input,    width = 23,                  .aruser
		.f2h_AWUSER           ()                                      //   input,    width = 23,                  .awuser
	);

	clk_100 clk_100 (
		.in_clk  (clk_100_clk),         //   input,  width = 1,  in_clk.clk
		.out_clk (clk_100_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	emif_calbus_0 emif_calbus_0 (
		.calbus_read_0          (emif_calbus_0_emif_calbus_0_calbus_read),    //  output,     width = 1,   emif_calbus_0.calbus_read
		.calbus_write_0         (emif_calbus_0_emif_calbus_0_calbus_write),   //  output,     width = 1,                .calbus_write
		.calbus_address_0       (emif_calbus_0_emif_calbus_0_calbus_address), //  output,    width = 20,                .calbus_address
		.calbus_wdata_0         (emif_calbus_0_emif_calbus_0_calbus_wdata),   //  output,    width = 32,                .calbus_wdata
		.calbus_rdata_0         (emif_hps_emif_calbus_calbus_rdata),          //   input,    width = 32,                .calbus_rdata
		.calbus_seq_param_tbl_0 (emif_hps_emif_calbus_calbus_seq_param_tbl),  //   input,  width = 4096,                .calbus_seq_param_tbl
		.calbus_clk             (emif_calbus_0_emif_calbus_clk_clk)           //  output,     width = 1, emif_calbus_clk.clk
	);

	emif_hps emif_hps (
		.pll_ref_clk          (emif_hps_pll_ref_clk_clk),                   //   input,     width = 1,     pll_ref_clk.clk
		.oct_rzqin            (emif_hps_oct_oct_rzqin),                     //   input,     width = 1,             oct.oct_rzqin
		.mem_ck               (emif_hps_mem_mem_ck),                        //  output,     width = 1,             mem.mem_ck
		.mem_ck_n             (emif_hps_mem_mem_ck_n),                      //  output,     width = 1,                .mem_ck_n
		.mem_a                (emif_hps_mem_mem_a),                         //  output,    width = 17,                .mem_a
		.mem_act_n            (emif_hps_mem_mem_act_n),                     //  output,     width = 1,                .mem_act_n
		.mem_ba               (emif_hps_mem_mem_ba),                        //  output,     width = 2,                .mem_ba
		.mem_bg               (emif_hps_mem_mem_bg),                        //  output,     width = 1,                .mem_bg
		.mem_cke              (emif_hps_mem_mem_cke),                       //  output,     width = 1,                .mem_cke
		.mem_cs_n             (emif_hps_mem_mem_cs_n),                      //  output,     width = 1,                .mem_cs_n
		.mem_odt              (emif_hps_mem_mem_odt),                       //  output,     width = 1,                .mem_odt
		.mem_reset_n          (emif_hps_mem_mem_reset_n),                   //  output,     width = 1,                .mem_reset_n
		.mem_par              (emif_hps_mem_mem_par),                       //  output,     width = 1,                .mem_par
		.mem_alert_n          (emif_hps_mem_mem_alert_n),                   //   input,     width = 1,                .mem_alert_n
		.mem_dqs              (emif_hps_mem_mem_dqs),                       //   inout,     width = 9,                .mem_dqs
		.mem_dqs_n            (emif_hps_mem_mem_dqs_n),                     //   inout,     width = 9,                .mem_dqs_n
		.mem_dq               (emif_hps_mem_mem_dq),                        //   inout,    width = 72,                .mem_dq
		.mem_dbi_n            (emif_hps_mem_mem_dbi_n),                     //   inout,     width = 9,                .mem_dbi_n
		.hps_to_emif          (agilex_hps_hps_emif_hps_to_emif),            //   input,  width = 4096,        hps_emif.hps_to_emif
		.emif_to_hps          (emif_hps_hps_emif_emif_to_hps),              //  output,  width = 4096,                .emif_to_hps
		.hps_to_emif_gp       (agilex_hps_hps_emif_gp_to_emif),             //   input,     width = 2,                .gp_to_emif
		.emif_to_hps_gp       (emif_hps_hps_emif_emif_to_gp),               //  output,     width = 1,                .emif_to_gp
		.calbus_read          (emif_calbus_0_emif_calbus_0_calbus_read),    //   input,     width = 1,     emif_calbus.calbus_read
		.calbus_write         (emif_calbus_0_emif_calbus_0_calbus_write),   //   input,     width = 1,                .calbus_write
		.calbus_address       (emif_calbus_0_emif_calbus_0_calbus_address), //   input,    width = 20,                .calbus_address
		.calbus_wdata         (emif_calbus_0_emif_calbus_0_calbus_wdata),   //   input,    width = 32,                .calbus_wdata
		.calbus_rdata         (emif_hps_emif_calbus_calbus_rdata),          //  output,    width = 32,                .calbus_rdata
		.calbus_seq_param_tbl (emif_hps_emif_calbus_calbus_seq_param_tbl),  //  output,  width = 4096,                .calbus_seq_param_tbl
		.calbus_clk           (emif_calbus_0_emif_calbus_clk_clk)           //   input,     width = 1, emif_calbus_clk.clk
	);

	qsys_top_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_100_out_clk_clk),                              //   input,   width = 1,   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //   input,  width = 10,     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //   input,   width = 1,       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //   input,   width = 1,       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //   input,   width = 1,       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //  output,  width = 32,       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //   input,  width = 32,       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //   input,   width = 4,       .byteenable
		.reset      (rst_controller_reset_out_reset),                   //   input,   width = 1, reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //   input,   width = 1,       .reset_req
	);

	qsys_top_pio_1 pio_1 (
		.clk        (clk_100_out_clk_clk),                   //   input,   width = 1,                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //   input,   width = 1,               reset.reset_n
		.address    (mm_interconnect_1_pio_1_s1_address),    //   input,   width = 2,                  s1.address
		.write_n    (~mm_interconnect_1_pio_1_s1_write),     //   input,   width = 1,                    .write_n
		.writedata  (mm_interconnect_1_pio_1_s1_writedata),  //   input,  width = 32,                    .writedata
		.chipselect (mm_interconnect_1_pio_1_s1_chipselect), //   input,   width = 1,                    .chipselect
		.readdata   (mm_interconnect_1_pio_1_s1_readdata),   //  output,  width = 32,                    .readdata
		.out_port   (fpga_led_pio_export)                    //  output,   width = 4, external_connection.export
	);

	rst_in rst_in (
		.clk         (clk_100_out_clk_clk),    //   input,  width = 1,       clk.clk
		.in_reset_n  (reset_reset_n),          //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (rst_in_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	user_rst_clkgate_0 user_rst_clkgate_0 (
		.ninit_done (ninit_done_ninit_done)  //  output,  width = 1, ninit_done.ninit_done
	);

	qsys_top_altera_mm_interconnect_1920_yigfcli mm_interconnect_0 (
		.agilex_hps_h2f_axi_master_awid                                             (agilex_hps_h2f_axi_master_awid),                   //   input,   width = 4,                                            agilex_hps_h2f_axi_master.awid
		.agilex_hps_h2f_axi_master_awaddr                                           (agilex_hps_h2f_axi_master_awaddr),                 //   input,  width = 32,                                                                     .awaddr
		.agilex_hps_h2f_axi_master_awlen                                            (agilex_hps_h2f_axi_master_awlen),                  //   input,   width = 8,                                                                     .awlen
		.agilex_hps_h2f_axi_master_awsize                                           (agilex_hps_h2f_axi_master_awsize),                 //   input,   width = 3,                                                                     .awsize
		.agilex_hps_h2f_axi_master_awburst                                          (agilex_hps_h2f_axi_master_awburst),                //   input,   width = 2,                                                                     .awburst
		.agilex_hps_h2f_axi_master_awlock                                           (agilex_hps_h2f_axi_master_awlock),                 //   input,   width = 1,                                                                     .awlock
		.agilex_hps_h2f_axi_master_awcache                                          (agilex_hps_h2f_axi_master_awcache),                //   input,   width = 4,                                                                     .awcache
		.agilex_hps_h2f_axi_master_awprot                                           (agilex_hps_h2f_axi_master_awprot),                 //   input,   width = 3,                                                                     .awprot
		.agilex_hps_h2f_axi_master_awvalid                                          (agilex_hps_h2f_axi_master_awvalid),                //   input,   width = 1,                                                                     .awvalid
		.agilex_hps_h2f_axi_master_awready                                          (agilex_hps_h2f_axi_master_awready),                //  output,   width = 1,                                                                     .awready
		.agilex_hps_h2f_axi_master_wdata                                            (agilex_hps_h2f_axi_master_wdata),                  //   input,  width = 32,                                                                     .wdata
		.agilex_hps_h2f_axi_master_wstrb                                            (agilex_hps_h2f_axi_master_wstrb),                  //   input,   width = 4,                                                                     .wstrb
		.agilex_hps_h2f_axi_master_wlast                                            (agilex_hps_h2f_axi_master_wlast),                  //   input,   width = 1,                                                                     .wlast
		.agilex_hps_h2f_axi_master_wvalid                                           (agilex_hps_h2f_axi_master_wvalid),                 //   input,   width = 1,                                                                     .wvalid
		.agilex_hps_h2f_axi_master_wready                                           (agilex_hps_h2f_axi_master_wready),                 //  output,   width = 1,                                                                     .wready
		.agilex_hps_h2f_axi_master_bid                                              (agilex_hps_h2f_axi_master_bid),                    //  output,   width = 4,                                                                     .bid
		.agilex_hps_h2f_axi_master_bresp                                            (agilex_hps_h2f_axi_master_bresp),                  //  output,   width = 2,                                                                     .bresp
		.agilex_hps_h2f_axi_master_bvalid                                           (agilex_hps_h2f_axi_master_bvalid),                 //  output,   width = 1,                                                                     .bvalid
		.agilex_hps_h2f_axi_master_bready                                           (agilex_hps_h2f_axi_master_bready),                 //   input,   width = 1,                                                                     .bready
		.agilex_hps_h2f_axi_master_arid                                             (agilex_hps_h2f_axi_master_arid),                   //   input,   width = 4,                                                                     .arid
		.agilex_hps_h2f_axi_master_araddr                                           (agilex_hps_h2f_axi_master_araddr),                 //   input,  width = 32,                                                                     .araddr
		.agilex_hps_h2f_axi_master_arlen                                            (agilex_hps_h2f_axi_master_arlen),                  //   input,   width = 8,                                                                     .arlen
		.agilex_hps_h2f_axi_master_arsize                                           (agilex_hps_h2f_axi_master_arsize),                 //   input,   width = 3,                                                                     .arsize
		.agilex_hps_h2f_axi_master_arburst                                          (agilex_hps_h2f_axi_master_arburst),                //   input,   width = 2,                                                                     .arburst
		.agilex_hps_h2f_axi_master_arlock                                           (agilex_hps_h2f_axi_master_arlock),                 //   input,   width = 1,                                                                     .arlock
		.agilex_hps_h2f_axi_master_arcache                                          (agilex_hps_h2f_axi_master_arcache),                //   input,   width = 4,                                                                     .arcache
		.agilex_hps_h2f_axi_master_arprot                                           (agilex_hps_h2f_axi_master_arprot),                 //   input,   width = 3,                                                                     .arprot
		.agilex_hps_h2f_axi_master_arvalid                                          (agilex_hps_h2f_axi_master_arvalid),                //   input,   width = 1,                                                                     .arvalid
		.agilex_hps_h2f_axi_master_arready                                          (agilex_hps_h2f_axi_master_arready),                //  output,   width = 1,                                                                     .arready
		.agilex_hps_h2f_axi_master_rid                                              (agilex_hps_h2f_axi_master_rid),                    //  output,   width = 4,                                                                     .rid
		.agilex_hps_h2f_axi_master_rdata                                            (agilex_hps_h2f_axi_master_rdata),                  //  output,  width = 32,                                                                     .rdata
		.agilex_hps_h2f_axi_master_rresp                                            (agilex_hps_h2f_axi_master_rresp),                  //  output,   width = 2,                                                                     .rresp
		.agilex_hps_h2f_axi_master_rlast                                            (agilex_hps_h2f_axi_master_rlast),                  //  output,   width = 1,                                                                     .rlast
		.agilex_hps_h2f_axi_master_rvalid                                           (agilex_hps_h2f_axi_master_rvalid),                 //  output,   width = 1,                                                                     .rvalid
		.agilex_hps_h2f_axi_master_rready                                           (agilex_hps_h2f_axi_master_rready),                 //   input,   width = 1,                                                                     .rready
		.onchip_memory2_0_s1_address                                                (mm_interconnect_0_onchip_memory2_0_s1_address),    //  output,  width = 10,                                                  onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                                  (mm_interconnect_0_onchip_memory2_0_s1_write),      //  output,   width = 1,                                                                     .write
		.onchip_memory2_0_s1_readdata                                               (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //   input,  width = 32,                                                                     .readdata
		.onchip_memory2_0_s1_writedata                                              (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //  output,  width = 32,                                                                     .writedata
		.onchip_memory2_0_s1_byteenable                                             (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //  output,   width = 4,                                                                     .byteenable
		.onchip_memory2_0_s1_chipselect                                             (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //  output,   width = 1,                                                                     .chipselect
		.onchip_memory2_0_s1_clken                                                  (mm_interconnect_0_onchip_memory2_0_s1_clken),      //  output,   width = 1,                                                                     .clken
		.agilex_hps_h2f_axi_reset_reset_bridge_in_reset_reset                       (~rst_in_out_reset_reset),                          //   input,   width = 1,                       agilex_hps_h2f_axi_reset_reset_bridge_in_reset.reset
		.agilex_hps_h2f_axi_master_translator_clk_reset_reset_bridge_in_reset_reset (~rst_in_out_reset_reset),                          //   input,   width = 1, agilex_hps_h2f_axi_master_translator_clk_reset_reset_bridge_in_reset.reset
		.clk_100_out_clk_clk                                                        (clk_100_out_clk_clk)                               //   input,   width = 1,                                                      clk_100_out_clk.clk
	);

	qsys_top_altera_mm_interconnect_1920_6idghsa mm_interconnect_1 (
		.agilex_hps_h2f_lw_axi_master_awid                                             (agilex_hps_h2f_lw_axi_master_awid),     //   input,   width = 4,                                            agilex_hps_h2f_lw_axi_master.awid
		.agilex_hps_h2f_lw_axi_master_awaddr                                           (agilex_hps_h2f_lw_axi_master_awaddr),   //   input,  width = 21,                                                                        .awaddr
		.agilex_hps_h2f_lw_axi_master_awlen                                            (agilex_hps_h2f_lw_axi_master_awlen),    //   input,   width = 8,                                                                        .awlen
		.agilex_hps_h2f_lw_axi_master_awsize                                           (agilex_hps_h2f_lw_axi_master_awsize),   //   input,   width = 3,                                                                        .awsize
		.agilex_hps_h2f_lw_axi_master_awburst                                          (agilex_hps_h2f_lw_axi_master_awburst),  //   input,   width = 2,                                                                        .awburst
		.agilex_hps_h2f_lw_axi_master_awlock                                           (agilex_hps_h2f_lw_axi_master_awlock),   //   input,   width = 1,                                                                        .awlock
		.agilex_hps_h2f_lw_axi_master_awcache                                          (agilex_hps_h2f_lw_axi_master_awcache),  //   input,   width = 4,                                                                        .awcache
		.agilex_hps_h2f_lw_axi_master_awprot                                           (agilex_hps_h2f_lw_axi_master_awprot),   //   input,   width = 3,                                                                        .awprot
		.agilex_hps_h2f_lw_axi_master_awvalid                                          (agilex_hps_h2f_lw_axi_master_awvalid),  //   input,   width = 1,                                                                        .awvalid
		.agilex_hps_h2f_lw_axi_master_awready                                          (agilex_hps_h2f_lw_axi_master_awready),  //  output,   width = 1,                                                                        .awready
		.agilex_hps_h2f_lw_axi_master_wdata                                            (agilex_hps_h2f_lw_axi_master_wdata),    //   input,  width = 32,                                                                        .wdata
		.agilex_hps_h2f_lw_axi_master_wstrb                                            (agilex_hps_h2f_lw_axi_master_wstrb),    //   input,   width = 4,                                                                        .wstrb
		.agilex_hps_h2f_lw_axi_master_wlast                                            (agilex_hps_h2f_lw_axi_master_wlast),    //   input,   width = 1,                                                                        .wlast
		.agilex_hps_h2f_lw_axi_master_wvalid                                           (agilex_hps_h2f_lw_axi_master_wvalid),   //   input,   width = 1,                                                                        .wvalid
		.agilex_hps_h2f_lw_axi_master_wready                                           (agilex_hps_h2f_lw_axi_master_wready),   //  output,   width = 1,                                                                        .wready
		.agilex_hps_h2f_lw_axi_master_bid                                              (agilex_hps_h2f_lw_axi_master_bid),      //  output,   width = 4,                                                                        .bid
		.agilex_hps_h2f_lw_axi_master_bresp                                            (agilex_hps_h2f_lw_axi_master_bresp),    //  output,   width = 2,                                                                        .bresp
		.agilex_hps_h2f_lw_axi_master_bvalid                                           (agilex_hps_h2f_lw_axi_master_bvalid),   //  output,   width = 1,                                                                        .bvalid
		.agilex_hps_h2f_lw_axi_master_bready                                           (agilex_hps_h2f_lw_axi_master_bready),   //   input,   width = 1,                                                                        .bready
		.agilex_hps_h2f_lw_axi_master_arid                                             (agilex_hps_h2f_lw_axi_master_arid),     //   input,   width = 4,                                                                        .arid
		.agilex_hps_h2f_lw_axi_master_araddr                                           (agilex_hps_h2f_lw_axi_master_araddr),   //   input,  width = 21,                                                                        .araddr
		.agilex_hps_h2f_lw_axi_master_arlen                                            (agilex_hps_h2f_lw_axi_master_arlen),    //   input,   width = 8,                                                                        .arlen
		.agilex_hps_h2f_lw_axi_master_arsize                                           (agilex_hps_h2f_lw_axi_master_arsize),   //   input,   width = 3,                                                                        .arsize
		.agilex_hps_h2f_lw_axi_master_arburst                                          (agilex_hps_h2f_lw_axi_master_arburst),  //   input,   width = 2,                                                                        .arburst
		.agilex_hps_h2f_lw_axi_master_arlock                                           (agilex_hps_h2f_lw_axi_master_arlock),   //   input,   width = 1,                                                                        .arlock
		.agilex_hps_h2f_lw_axi_master_arcache                                          (agilex_hps_h2f_lw_axi_master_arcache),  //   input,   width = 4,                                                                        .arcache
		.agilex_hps_h2f_lw_axi_master_arprot                                           (agilex_hps_h2f_lw_axi_master_arprot),   //   input,   width = 3,                                                                        .arprot
		.agilex_hps_h2f_lw_axi_master_arvalid                                          (agilex_hps_h2f_lw_axi_master_arvalid),  //   input,   width = 1,                                                                        .arvalid
		.agilex_hps_h2f_lw_axi_master_arready                                          (agilex_hps_h2f_lw_axi_master_arready),  //  output,   width = 1,                                                                        .arready
		.agilex_hps_h2f_lw_axi_master_rid                                              (agilex_hps_h2f_lw_axi_master_rid),      //  output,   width = 4,                                                                        .rid
		.agilex_hps_h2f_lw_axi_master_rdata                                            (agilex_hps_h2f_lw_axi_master_rdata),    //  output,  width = 32,                                                                        .rdata
		.agilex_hps_h2f_lw_axi_master_rresp                                            (agilex_hps_h2f_lw_axi_master_rresp),    //  output,   width = 2,                                                                        .rresp
		.agilex_hps_h2f_lw_axi_master_rlast                                            (agilex_hps_h2f_lw_axi_master_rlast),    //  output,   width = 1,                                                                        .rlast
		.agilex_hps_h2f_lw_axi_master_rvalid                                           (agilex_hps_h2f_lw_axi_master_rvalid),   //  output,   width = 1,                                                                        .rvalid
		.agilex_hps_h2f_lw_axi_master_rready                                           (agilex_hps_h2f_lw_axi_master_rready),   //   input,   width = 1,                                                                        .rready
		.pio_1_s1_address                                                              (mm_interconnect_1_pio_1_s1_address),    //  output,   width = 2,                                                                pio_1_s1.address
		.pio_1_s1_write                                                                (mm_interconnect_1_pio_1_s1_write),      //  output,   width = 1,                                                                        .write
		.pio_1_s1_readdata                                                             (mm_interconnect_1_pio_1_s1_readdata),   //   input,  width = 32,                                                                        .readdata
		.pio_1_s1_writedata                                                            (mm_interconnect_1_pio_1_s1_writedata),  //  output,  width = 32,                                                                        .writedata
		.pio_1_s1_chipselect                                                           (mm_interconnect_1_pio_1_s1_chipselect), //  output,   width = 1,                                                                        .chipselect
		.agilex_hps_h2f_lw_axi_reset_reset_bridge_in_reset_reset                       (~rst_in_out_reset_reset),               //   input,   width = 1,                       agilex_hps_h2f_lw_axi_reset_reset_bridge_in_reset.reset
		.agilex_hps_h2f_lw_axi_master_translator_clk_reset_reset_bridge_in_reset_reset (~rst_in_out_reset_reset),               //   input,   width = 1, agilex_hps_h2f_lw_axi_master_translator_clk_reset_reset_bridge_in_reset.reset
		.clk_100_out_clk_clk                                                           (clk_100_out_clk_clk)                    //   input,   width = 1,                                                         clk_100_out_clk.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~rst_in_out_reset_reset),            //   input,  width = 1, reset_in0.reset
		.clk            (clk_100_out_clk_clk),                //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //  output,  width = 1,          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

endmodule
